library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is 
	port(
		cord_x    : in std_logic_vector (2 downto 0);
		cord_y    : in std_logic_vector (2 downto 0);
		digito: in std_logic_vector (3 downto 0);
		rom_out       : out std_logic
		);
end;

architecture ROM_arq of ROM is
type matriz is array (0 to 95) of std_logic_vector(0 to 7);
	signal direc: std_logic_vector(6 downto 0);
	
constant caracteres: matriz :=("00000000",
							   "00111100", 
							   "01000010", 
							   "01000010", 
							   "01000010", 
							   "01000010", 
							   "00111100", 
							   "00000000", 	--0

							   "00000000",
							   "00001000",
							   "00011000",
						       "00001000",
							   "00001000",
							   "00001000",
							   "00001000",
							   "00000000", --1

							   "00000000",
							   "00111100",
							   "01000010",
							   "00000100",
							   "00001000",
							   "00110000",
							   "01111110",
							   "00000000", --2

							   "00000000",
						       "01111100",
							   "00000010",
							   "00111100",
							   "00000010",
							   "00000010",
							   "01111100",
							   "00000000",--3

							   "00000000",
							   "00001100",
							   "00010100",
							   "00100100",
							   "01111110",
							   "00000100",
							   "00000100",
							   "00000000",--4

							   "00000000",
							   "01111110",
							   "01000000",
							   "01111100",
							   "00000010",
							   "00000010",
							   "01111100",
							   "00000000",--5

							   "00000000",
							   "00111110",
							   "01000000",
							   "01111100",
							   "01000010",
							   "01000010",
							   "00111100",
							   "00000000",--6

							   "00000000",
							   "01111110",
							   "00000110",
							   "00001000",
							   "00010000",
							   "00100000",
							   "00100000",
							   "00000000",--7

							   "00000000",
							   "00111100",
							   "01000010",
							   "00111100",
							   "01000010",
							   "01000010",
							   "00111100",
							   "00000000",--8

							   "00000000",
							   "00111100",
							   "01000010",
							   "01000010",
							   "00111110",
							   "00000010",
							   "00011100",
							   "00000000",--9

							   "00000000",
							   "00000000",
							   "00000000",
							   "00000000",
							   "00000000",
							   "00011000",
							   "00011000",
							   "00000000",--.

							    "00000000", 
								"01000010", 
								"01100110", 
								"01100110", 
							    "01100110", 
								"00111100", 
								"00011000", 
								"00000000");--V
								
begin
	direc  <= digito & cord_x;	
	rom_out  <= caracteres(to_integer(unsigned(direc)))(to_integer(unsigned(cord_y)));

end;